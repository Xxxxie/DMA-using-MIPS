LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY MUX31 IS
PORT ( 
 Rs  : IN  STD_LOGIC_VECTOR(4 DOWNTO 0 );
  Rt  : IN  STD_LOGIC_VECTOR(4 DOWNTO 0 );
  Rd  : IN  STD_LOGIC_VECTOR(4 DOWNTO 0 ); 
T1,T2 : IN STD_LOGIC;
isRead : IN STD_LOGIC;
COUT : OUT STD_LOGIC_VECTOR(4 DOWNTO 0)

 );
END MUX31;
ARCHITECTURE behav OF MUX31 IS

BEGIN

PROCESS(Rs,Rt,Rd,T1,T2,isRead)
BEGIN

if T1='1' then COUT<=Rs; 
else if T2='1'then COUT<=Rt; 
 else  COUT<=Rd;  
end if;
end if;

END PROCESS;

END behav;
