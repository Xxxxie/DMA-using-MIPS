LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY ALU IS
PORT ( S  : IN  STD_LOGIC_VECTOR(5 DOWNTO 0 );
A,B  : IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
F  : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
Z : OUT STD_LOGIC;
CN  : IN  STD_LOGIC
  );
END ALU;
ARCHITECTURE behav OF ALU IS
SIGNAL A32,B32,F32 : STD_LOGIC_VECTOR(31 DOWNTO 0);
BEGIN

PROCESS(CN,A32,B32)
BEGIN
Z <='1';
CASE S  IS
WHEN "000000" => F32<=A32;
WHEN "000010" => F32<=A + B+ CN; 
WHEN "000110" => F32<= A - B;
				if (F32 = "00000000000000000000000000000000") then Z <='0';
				END IF;
WHEN "000011" => F32<=A and B;
WHEN "000001" => F32<=A or B;              
WHEN OTHERS  =>F32<= "00000000000000000000000000000000" ;
END CASE;

END PROCESS;
F<= F32(31 DOWNTO 0) ;  

END behav;
